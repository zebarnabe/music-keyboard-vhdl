----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:10:16 07/01/2015 
-- Design Name: 
-- Module Name:    keyMatrixLED - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity keyMatrixLED is
    Port ( keyMatrix : in  STD_LOGIC_VECTOR (31 downto 0);
           led : out  STD_LOGIC_VECTOR (7 downto 0));
end keyMatrixLED;

architecture Behavioral of keyMatrixLED is
begin
  led <= (keyMatrix(31 downto 24) xor keyMatrix(23 downto 16) xor keyMatrix(15 downto 8) xor keyMatrix(7 downto 0));
end Behavioral;

